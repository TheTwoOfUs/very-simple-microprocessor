CIRCUIT D:\Documents and Settings\sicard\Mes documents\microwind31\examples\AmpliFollow.MSK
*
* IC Technology: CMOS 0.12�m - 6 Metal
*
VDD 1 0 DC 1.20
VV+ 9 0 DC 0 PULSE(0.38 0.67 4.10N 0.10N 0.10N 4.10N 8.40N)
*
* List of nodes
* "out" corresponds to n�3
* "N4" corresponds to n�4
* "N5" corresponds to n�5
* "N6" corresponds to n�6
* "N8" corresponds to n�8
* "V+" corresponds to n�9
* "Vref" corresponds to n�10
*
* MOS devices
MN1 0 5 5 0 N1  W= 0.36U L= 0.12U
MN2 3 5 0 0 N1  W= 0.36U L= 0.12U
MN3 8 9 4 0 N1  W= 0.36U L= 0.12U
MN4 0 1 8 0 N1  W= 1.08U L= 0.12U
MN5 6 3 8 0 N1  W= 0.36U L= 0.12U
MP1 1 4 3 1 P1  W= 0.84U L= 0.12U
MP2 4 4 1 1 P1  W= 0.84U L= 0.12U
MP3 1 6 5 1 P1  W= 0.84U L= 0.12U
MP4 6 6 1 1 P1  W= 0.84U L= 0.12U
*
C2 1 0  4.182fF
C3 3 0  1.260fF
C4 4 0  0.745fF
C5 5 0  1.152fF
C6 6 0  0.692fF
C8 8 0  0.519fF
C9 9 0  0.171fF
C10 1 0  0.145fF
*
* Extra RLC
*
Cadd1 3 0 1pF
*
*
* n-MOS BSIM4 :
* low leakage
.MODEL N1 NMOS LEVEL=14 VTHO=0.40 U0=0.050 TOXE= 2.0E-9 LINT=0.010U 
+K1 =0.450 K2=0.100 DVT0=2.300
+DVT1=0.540 LPE0=23.000e-9 ETA0=0.080
+NFACTOR=  1.6 U0=0.050 UA=3.000e-15
+WINT=0.020U LPE0=23.000e-9 
+KT1=-0.060 UTE=-1.800 VOFF=0.050
+XJ=0.150U NDEP=170.000e15 PCLM=1.100
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p
*
* p-MOS BSIM4:
* low leakage
.MODEL P1 PMOS LEVEL=14 VTHO=-0.45 U0=0.018 TOXE= 2.0E-9 LINT=0.010U 
+K1 =0.450 K2=0.100 DVT0=2.300
+DVT1=0.540 LPE0=23.000e-9 ETA0=0.080
+NFACTOR=  1.6 U0=0.018 UA=1.500e-15
+WINT=0.020U LPE0=23.000e-9 
+KT1=-0.060 UTE=-1.800 VOFF=0.050
+XJ=0.150U NDEP=170.000e15 PCLM=0.700
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p
*
* Transient analysis
*
* (Winspice)
.options temp=27.0
.control
tran 0.1N 20.00N
print  V(9) V(3) > out.txt
plot  V(9) V(3)
.endc
.END
